module serialAdder_tb();
    
endmodule