module serialAdder ();

// pg. 653 on the txtbook
    
endmodule