module top();
    
endmodule