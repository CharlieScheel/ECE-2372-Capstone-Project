module top;

/* declare variables here */
reg zFlag,      // Equals 1 if the result of the subtraction operation is 0x00
    nFlag,      // Equals 1 if the result of the subtraction is negative
    vFlag;      // Equals 1 if the subtraction operation results in an overflow
reg [7:0] a;    // Accumulator
reg [7:0] b;    // Subtrahend register

initial begin
    
    /*

    */

end

endmodule


module serialAdder ();

// pg. 653 on the txtbook
    
endmodule


module top_tb();
    
endmodule


module serialAdder_tb();
    
endmodule